module DM(
	input clk,
	input WE,
	input [31:0] A,
	input [31:0] WD,
	output [31:0] RD
);